module Text;
    initial $display("Hello World!");
endmodule